module main

import time

fn hello() string {
	return 'Hello world'
}

fn main() {
	hello()
}
